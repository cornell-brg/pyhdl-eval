//========================================================================
// const_ref
//========================================================================
// SPDX-License-Identifier: MIT
// Author : Christopher Batten, NVIDIA
// Date   : May 20, 2024

module RefModule
(
  output logic [7:0] out
);

  assign out = 1;

endmodule

